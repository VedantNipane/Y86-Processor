`timescale 1ns / 1ps

module not1x1(
  input  a,
  output  out
  );

  not gate1(out,a);  

endmodule