`timescale 1ns / 1ps

module and1x1(
  input  a,
  input  b,
  output  out
  );

  and g1(out,a,b);  

endmodule